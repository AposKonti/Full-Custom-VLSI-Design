* File: /home/eng/a/axk220238/vlsi/cad/gf65/axk220238_axk230133/AOI22/AOI22_lvs/AOI22.pex.sp
* Created: Thu Nov 30 17:45:52 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "AOI22.pex.sp.pex"
.subckt AOI22  VSS OUT VDD IN1 IN2 IN3 IN4
* 
* IN4	IN4
* IN3	IN3
* IN2	IN2
* IN1	IN1
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=4.43025e-12
+ PERIM=8.53e-06
XMMN0 NET17 N_IN1_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.2e-07 AD=5.2e-14 AS=8.788e-14 PD=7.2e-07 PS=1.378e-06 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.69e-07
+ SB=9.55e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMN1 N_OUT_MMN1_d N_IN2_MMN1_g NET17 N_VSS_D0_noxref_pos NFET L=6.4e-08
+ W=5.2e-07 AD=5.226e-14 AS=5.2e-14 PD=7.21e-07 PS=7.2e-07 NRD=0.194231
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=4.34e-07
+ SB=6.91e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.6e-15 PANW4=3.2e-15 PANW5=3.2e-15
+ PANW6=6.4e-15 PANW7=1.28e-14 PANW8=6.08e-15 PANW9=0 PANW10=0
XMMN2 N_OUT_MMN1_d N_IN3_MMN2_g NET026 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.2e-07 AD=5.226e-14 AS=5.2e-14 PD=7.21e-07 PS=7.2e-07 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=6.99e-07
+ SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMN3 NET026 N_IN4_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.2e-07 AD=5.2e-14 AS=8.32e-14 PD=7.2e-07 PS=1.36e-06 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=9.64e-07
+ SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMP0 N_NET11_MMP0_d N_IN1_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=1.5548e-13 AS=9.2e-14 PD=2.178e-06 PS=1.12e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.69e-07 SB=9.55e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.63e-14 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=9.3275e-14
+ PANW10=3.9e-14
XMMP1 N_NET11_MMP1_d N_IN2_MMP1_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=9.2e-14 PD=1.12e-06 PS=1.12e-06 NRD=0.108696
+ NRS=0.108696 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1 SA=4.34e-07
+ SB=6.9e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=2.588e-14 PANW8=1.1604e-13 PANW9=3.7155e-14 PANW10=3.9e-14
XMMP2 N_OUT_MMP2_d N_IN3_MMP2_g N_NET11_MMP1_d N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=9.2e-14 PD=1.12e-06 PS=1.12e-06 NRD=0.108696
+ NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=6.99e-07
+ SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=7.28e-14 PANW8=1.3e-14 PANW9=9.3275e-14 PANW10=3.9e-14
XMMP3 N_OUT_MMP2_d N_IN4_MMP3_g N_NET11_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=1.472e-13 PD=1.12e-06 PS=2.16e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=9.64e-07 SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=4.097e-14
+ PANW5=2.533e-14 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=9.3275e-14
+ PANW10=3.9e-14
c_156 NET026 0 3.50179e-20
*
.include "AOI22.pex.sp.AOI22.pxi"
*
.ends
*
*

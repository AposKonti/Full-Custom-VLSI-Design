* File: /home/eng/a/axk220238/vlsi/cad/gf65/axk220238_axk230133/NAND/NAND_lvs/NAND.pex.sp
* Created: Thu Nov 30 17:59:12 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "NAND.pex.sp.pex"
.subckt NAND  VSS OUT VDD IN1 IN2
* 
* IN2	IN2
* IN1	IN1
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=2.81655e-12
+ PERIM=7.226e-06
XMMN0 NET15 N_IN1_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.2e-07 AD=5.2e-14 AS=8.32e-14 PD=7.2e-07 PS=1.36e-06 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.6e-07
+ SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMN1 N_OUT_MMN1_d N_IN2_MMN1_g NET15 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.2e-07 AD=8.32e-14 AS=5.2e-14 PD=1.36e-06 PS=7.2e-07 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.25e-07
+ SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMP0 N_OUT_MMP0_d N_IN1_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=1.472e-13 PD=1.12e-06 PS=2.16e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.6e-07 SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=4.557e-14
+ PANW5=2.073e-14 PANW6=6.5e-15 PANW7=7.28e-14 PANW8=1.3e-14 PANW9=3.3475e-14
+ PANW10=3.9e-14
XMMP1 N_OUT_MMP0_d N_IN2_MMP1_g N_VDD_MMP1_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=1.472e-13 PD=1.12e-06 PS=2.16e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=4.25e-07 SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=4.557e-14
+ PANW5=2.073e-14 PANW6=6.5e-15 PANW7=7.28e-14 PANW8=1.3e-14 PANW9=3.3475e-14
+ PANW10=3.9e-14
c_42 NET15 0 3.48696e-20
*
.include "NAND.pex.sp.NAND.pxi"
*
.ends
*
*

* File: /home/eng/a/axk220238/vlsi/cad/gf65/axk220238_axk230133/OR/OR_lvs/OR.pex.sp
* Created: Thu Nov 30 18:08:58 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "OR.pex.sp.pex"
.subckt OR  OUT VSS VDD IN1 IN2
* 
* IN2	IN2
* IN1	IN1
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=3.6531e-12
+ PERIM=7.902e-06
XMMN3 N_OUT_MMN3_d N_NET07_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.2e-07 AD=8.32e-14 AS=5.2e-14 PD=1.36e-06 PS=7.2e-07 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.6e-07
+ SB=6.9e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMN0 N_NET07_MMN0_d N_IN1_MMN0_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.2e-07 AD=5.2e-14 AS=5.2e-14 PD=7.2e-07 PS=7.2e-07 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=4.25e-07
+ SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMN1 N_NET07_MMN0_d N_IN2_MMN1_g N_VSS_MMN1_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.2e-07 AD=5.2e-14 AS=8.32e-14 PD=7.2e-07 PS=1.36e-06 NRD=0.192308
+ NRS=0.192308 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=6.9e-07
+ SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=6.175e-15 PANW9=0 PANW10=0
XMMP3 N_OUT_MMP3_d N_NET07_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=1.472e-13 AS=9.2e-14 PD=2.16e-06 PS=1.12e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.6e-07 SB=6.9e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15
+ PANW5=2.441e-14 PANW6=4.514e-14 PANW7=1.3e-14 PANW8=7.28e-14 PANW9=3.3475e-14
+ PANW10=3.9e-14
XMMP0 N_NET012_MMP0_d N_IN1_MMP0_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=9.2e-14 AS=9.2e-14 PD=1.12e-06 PS=1.12e-06 NRD=0.108696
+ NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=4.25e-07
+ SB=4.25e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.2616e-13 PANW8=1.944e-14 PANW9=3.3475e-14 PANW10=3.9e-14
XMMP1 N_NET07_MMP1_d N_IN2_MMP1_g N_NET012_MMP0_d N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.2e-07 AD=1.472e-13 AS=9.2e-14 PD=2.16e-06 PS=1.12e-06
+ NRD=0.108696 NRS=0.108696 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1
+ SA=6.9e-07 SB=1.6e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.625e-15 PANW4=4.557e-14
+ PANW5=2.073e-14 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=9.3275e-14
+ PANW10=3.9e-14
*
.include "OR.pex.sp.OR.pxi"
*
.ends
*
*
